module datapath
	(
		input resetn,
		input clk,
		input [3:0] keypress,
		input [3:0] songselect,
		input initialize,
		input ld_notes,
		input erase_notes,
		input draw_board,
		input draw_notes1,
		input draw_notes2,
		input draw_notes3,
		input draw_notes4,
		input check_notes,
		input playerEN,
		input [3:0] song,
		output reg [818:0] song_note1,
		output reg [818:0] song_note2,
		output reg [818:0] song_note3,
		output reg [818:0] song_note4,
		output reg [7:0] x_out,
		output reg [7:0] y_out,
		output reg [2:0] colour_out,
		output reg [15:0] score,
		output reg done,
		output reg updating
	);
			
	
	reg [7:0] x_coordinate;
	reg [7:0] y_coordinate;
	
	reg [119:0] note1_bar;
	reg [119:0] note2_bar;
	reg [119:0] note3_bar;
	reg [119:0] note4_bar;
	reg [17:0] counter;
	reg [7:0] offset;
	
	reg [2:0] shift_counter;
	reg [7:0] x_board_counter;
	reg [7:0] y_board_counter;
	reg [3:0] line_counter;
	
	reg [3:0] next_note;
	reg [3:0] hold_note;
	
	reg [7:0] temp_score1;
	reg [7:0] temp_score2;
	reg [7:0] temp_score3;
	reg [7:0] temp_score4;
	
	always @(posedge clk)
	begin
		if(!resetn)
		begin
			colour_out <= 3'b000;
			offset <= 8'b0;
			counter <= 8'b0;
			note1_bar <= 120'b0;
			note2_bar <= 120'b0;
			note3_bar <= 120'b0;
			note4_bar <= 120'b0;
			done <= 1'b0;
			updating <= 1'b0;
			
			if(counter < 17'b1000_0000_0000_0000_0)
			begin
				counter <= counter + 1'b1;
				x_coordinate <= counter[7:0];
				y_coordinate <= counter[15:8];
			end
			else
			begin
				counter <= 0;
				x_coordinate <= 8'b0;
				y_coordinate <= 8'b0;
			end
				
		end
		
		if(initialize)
		begin
			score <= 8'b0;
			shift_counter <= 3'b000;
			temp_score1 <= 8'b0;
			temp_score2 <= 8'b0;
			temp_score3 <= 8'b0;
			temp_score4 <= 8'b0;
			
			x_coordinate <= 8'b0;
			y_coordinate <= 8'b0;
			
			if(song == 4'b0001)
			begin
				song_note1 <= 819'b1001001001001001001001000000000000001000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001000000000000001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010000000001001001001001001001001001001001001001001001001000100010010100001001001001000000000000001001001001000000000001000000000001000000000000000000000000000000000000100010101001111110100101111110100101111110100101001001001001000000001000100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100100000000000100100100100100000000000000000001001100000000000000000001100100001010001010001000000000001111110111111111111;
				song_note2 <= 819'b0100100100100100100100101001001001000100100100100100100100010100100100010100100100010100100100010100100100010100100100010100100100010100100100010100100100011001001001000100100100010100100100010100100100010100100100010100100100010100100100010100100100010100100100010000101000000100100100010100100100010100100100010100100100010010001000010100100100100100100100101000100100010010101000010010101000010010101000011000101000100100010100010010100010100100100100100100100100100100100100100100100100100101001000100010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010100100100010010010010010010100001100001010100101010100001100010100001010010001010001010000000000001111110111111111111;
				song_note3 <= 819'b0010010010010010010010010100100100100010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010100100100010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010010000000010100010010010010010010010010010010010010010010010010001000100000010010010010010010010010100000010000101000010100101000010010101000010010010100100100010100010101000101000010010100001010010100001010010100001010010010010010010100100010001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001001010010010001001001001001010001010001010100100010100001010001001010010100100000100000100000000000001111110111111111111;
				song_note4 <= 819'b0000000000000000000000000010010010010001000001111111111101011111101111111111101001001000000000000000000001011111110001011111110000011111110001011111110111110010010010011111111110101111111110101111111110101111101111111111101111111111101111111111101111111111110010100000000000001111110001011111110010101111111110101111110010101000000001010000000000000001001001000000010000000000010100010000010100100000010100010100010100011000101000100000000000000000000000000000000000000000000000000000000000000000010010111111111110101111110111111111110100100100000001001111111101001111110001001111110111111011110111111011111100100011111100100011111100100011111100100111110111110011111110100100100100100111110100100100001001001000000000000000001010100010100010010000001010100010100000000000000000000000000000000000000000000000000000000;
			end
			else if(song == 4'b0010)
			begin
				song_note1 <= 819'b1001011110100110010100010010110101010011011111011011110000011110011000100111000010110001110011101011010000011011110111101100001011110100111101111110110110110001110010101101001110010101010100000000110101011000111110011101100010010010110011111111000110010000001111011001101101011110000110110011010100001100001100011100100101111010000011001100101010010001011110000010011110101100100010101110011011000100000010001010001010110001111110010100101000110101000011110101111100100110110011011001111001100011000000111000000101001110100011000110011110000111001110010010101101101101011111000110001011010011001100010010110110110010000101010011110100010001111100001010000011010000011100101010111011001110110000110010010111100011010100110110011101010111000010111001100100111100110101111100111000111001100101001101110110001101000010001;
				song_note2 <= 819'b1111101101011011000001010001111110110101111101110011011100000001100100100010011110101011000111111010100101111100010010011111011001010100001010001000101110010001100011000100110101011110110000101111111011100010110000010100011000110101111111011011101010110100110010110000110100101111010000110110111011001010010000101010010100000110100011111111101110001101001010011000111100101011010100100100000110001000100110011111001001110111010110001100101010011011111010011010000010100000010000001011100000001001000001111000101100101001111011100101100110001100010100111110001101010000110011101011110101000100101100100000011110110110010110111111000111011000110110100110011101010001001101100101100000100011111000001001100000101010000000010010111101010001100000100100010111111101001100011100010110100111110100001011011010011100110000011;
				song_note3 <= 819'b0010111010101010101011011000111010010100001000100011101000110100111111110101101001011000110010000110001111001011001000011011000011010000000111000111000001010111101010000100111111100001011111010000001111100111110011111110000011100110100101000100010101110110000000011111101010110111000110100000100101111010010100101100011101100110001110110000110010000110000000001100100110100101010111111111111101101011010001001001000000111101011100111111010000000011011111111011101001101111010111011011100010011011101100101001011000110100111110111001100101110001011111110000110111010110010001011101110000111110111100111000011110111111101000100100000000111010101001100111001100011101100100001011101111111011100010010111000011110101100101000001110101001001111101010010011111101010011110010110101111001001011010110010101011111010101010111;
				song_note4 <= 819'b0101010011011111111000010010010010010101110000101000001001100101101011101011010000100111111100000101101101111111101101111111101110011111001001100111001111011010101010101000001101101110001111111011100100101101110100010110011111110101011000001011001000001011101000111001010001110010000101100000110011011111010010011100101111011111111111100010101101100111101010001100101101001010010110110011100110111011001010100010100010111001100110100010011111001111010011011100101001001100010110010011011010000001001111110110111101101011111101010000110001101101100000000010011000001011111000101010110001011110101010100111010011111101010101101111100101011101100010101001111001111100001001111100000001010000110011110011000010010111011011101110000100101011010100101100101011000101100111000011000110111001010111111000001101110101011000011;
			end
			else if(song == 4'b0011)
			begin
				song_note1 <= 819'b0001000000000010000000001000000000000001000010110001000001010000000000000000100000000000011010000001000010001000000000000000000010000100000001000101000000010000001000101000010100000000100010001000010001000010001111010100000000000001011011010000001000100010000000100000000011100100100110111000100000011010100001000000000100011001000000010000000010101011000010100010000000000000000001001101100000000000000100000111011000001000000000010100001000011010000001001001000100010000010000000000000000001110000001001110000000000000011010000001010000000001101100000100011010101100101110011000100010000001000110000011000000010000011000000000000110000000010001000000000001010000011010001110000000100101000000000110000101000011000000100000011110011001101000100000000000001011001000000001100000001110100000000010000001000011100000100;
				song_note2 <= 819'b0001000000010001001000000001000000000010101010000000001010000110100001000000110000001000000000000000000010100001000000000011000010000001100110010010000000000001001001010100001000000000000000000000000001000000000001000100000000101011001000010000100110000110010000000000000000000000000001000000000010100100000000001000000101000000100000000001000100001000000000000000110000100000100010000110011000000000000011000000000000100000101000011100110000000001000000110000000000000000000000001100010001010000010000000001000000100010000000010010010010000000000000000000000100000000010000010000000000010100100001000000000001000010000000000000100110000100000100100000000100000010000010001000000000001100010000000000000000000000001001010010000000000000000100001000000000000010100000001000000001101010100001000000000111000001001000000;
				song_note3 <= 819'b0000000001000000000000010000010000100100000000000000111100000000000000000000100000001010000000100101100001011010110101101000100001000010000010011010000001000000000010100101000101010000010011000000000000010000000000000001000010110000000000001000100100010000000000011000000000010000001100000001000010000010000111001100000000000001011111100100100000000010000000000000101100100001000010100000000000000000000100100011000000001000000100110000100000001000100001000000010000111100000000000001000000000001110000000100011000100000010001000000010000000011000000001000001100000100010000010000000000001000010010010101010000000001000100000001000111010000000001011000000100001000000000010111000000000010010101110010010010010010000000000000000000000000000000011101001100010001101010010000000000101000000000000001001010100011000000010;
				song_note4 <= 819'b0000110000000000110100100001000010000010000000001110000001000001100000000000100000101000001000000000000001010000110000000001000000000100000000000000000000100010001000000000000110000000000010000100000000000101000000001001000100100000000100001000001000001000000100010000101000010000101000100010000000000001010010000000000010011000000000000000001111011001000100000100001000000011001000001000110000101010100010000100000100000000010000011000100001100001000001000000000010000001000000000110100000000100000000001001010000011010010001100100001101000011010010001010000000001000000000000000001000001000111000001000001110100000000000100000000011001000000010000001000000001010000010001000001000001001010100000100010110000000000001000000000100000000000000111010000110101000010001100010010010100010000010100101000100000000001000100;
			end
			else if(song == 4'b0100)
			begin
				song_note1 <= 819'b0000000000000000010100000000000100000001000000000000000000010000000010100000000000000000000001000000000000010000000001000000000010000000000000000000000000001000001000000100100000000000000000000000000000100000000000000000000001010000000000000000000000000000000000000000000000000000000000100000000000001000000010000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000100000000000000010000000000000000000000100100000000000000000000000000000000000100000000000000000001000000000000000001000100000000000000000000010100001000000000000000000000000000000000010100000000000000000000000000000000000100000000001000000000000000000000000000000000000000100000000000000000000000000000000000001000100000000000000000000000001000001000010000010000000000000000001010000000000000000000000000000000001000;
				song_note2 <= 819'b0000100000000000000000000000100000000000010000000000000000000001010000000000010000000000000000000000010000001000011000010000000000001000000001000000000000000000000000000000000000000100000000000000000000000000000000000100001000000100000000000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000000100000010000000000000000100000000000000000000000000100000100000000000000000000000000000010000000000000000010000000000000000001000000000110000000000000000000000000000000000000001000000010100100000000000000000000000000000000000001000000000000000000000000000000100000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000100100010000000000000000000000000001000000000000000100000000000100000000000010001000000000000000000000001000000000;
				song_note3 <= 819'b0000000000000000000000000000000100000100000000001000010001000000000000000001000000000000000100000000000000000001000000000000100000000000000000000000000010000000000000000000010000000000000001000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000011000000010000000000000010010000000000000000000000000000000000000010000000000000001100001000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000010000000000000000000000000000000100000000010000000000000000000010000000000010100000000000000000000110000100000000000000100000000000000100000000000000000000000000000000000000000000010000000000001000000100000000000100000001000000000000000000000000000010000001000000000100000000001;
				song_note4 <= 819'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000100101100000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000010000000000000000000100000000000100000000000000100010000000000000000000000000000010000000000000000000000000000100000000000000000001000000000000010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000001000000000100100000000100000000000000100000000000000000001000000000000000000000000000000010000000000000000000000001000100000000000000;
			end
			else if(song == 4'b0101)
			begin
				song_note1 <= 819'b0000000100000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000100000001010000000000000000000000000000000000000000000000000000000010000000000010000000000000000000000000000000000100010000000000000000010000000000000001000000000000000000000000000000100000000100000000000000000011000000000000000000000000000001000000000000100000000010000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000001000000000000000000000000000000000000000000000000000000001000;
				song_note2 <= 819'b0000000000000000000100000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000010000000000000000000000000000000000000000000000010010000000000000000000000000000010000000000000000000000000000000000000000000001000000000000000000000000000000001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000100000001000000000000000000000000100000000000000000000000000100000000000000010000000100000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000100001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000;
				song_note3 <= 819'b0000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000010000000000000000000000000000000000000000000100000000000100000000000000000000000000000000001000000000000000000000000001000000010000000000000000000000000000000000000100000000000000000000000000000000100001000000000000000000000000000000000100000000000000100000;
				song_note4 <= 819'b0000000000000000000000000000000000000000000100000000000000100001010000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000100000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000100000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000100000000000000000000000000000001000000000000000000000001000000000000000000010000000000000000000000000000000000000000000000000000000000000000000;
			end
			else if(song == 4'b0110)
			begin
				song_note1 <= 819'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000000000000000000000000000010010000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000010000000000000000000000000000000000000010001000000000000000000000000100000000000000000000000000000000000001000;
				song_note2 <= 819'b0000000000000000000000000000000000000000000000000000000000000000000100000000001000010000000000000100000000000000000000000000000000000000000000000000000000000100000000000000000000000000010000000001000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100011000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
				song_note3 <= 819'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000001000000000000000000000000000000000000000000000000000010010100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000100001100000000000000000000000000000000000000010000000000001000000000000000000000000000010000000000000000000000000000000000000000000010000000000001000000000000000000010000000000000000000000000000101000000000000000000000000000000000000000000001000000000000000000010000000000;
				song_note4 <= 819'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000000000000000010010000000000000000000000000000000000000000000000100000000000010000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000100000000000000000000000000001000000000000000000000000000000000000000000000000000000000000100001000000000000000000000000000000000000010000000000100000000000;
			end
			else if(song == 4'b0111)
			begin
				song_note1 <= 819'b0000000000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000010010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000010000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				song_note2 <= 819'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
				song_note3 <= 819'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000100000000000000000000000000000000000000000000000000;
				song_note4 <= 819'b0000000010000000000000000000000000000000001000000000000000000000001000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			end
			else
			begin
				song_note1 <= 819'b0;
				song_note2 <= 819'b0;
				song_note3 <= 819'b0;
				song_note4 <= 819'b0;
			end
			
		end
			
		if(ld_notes)
		begin
		
			line_counter <= 4'b0000;
			colour_out <= 3'b000;
			x_coordinate <= 8'b0;
			y_coordinate <= 8'b0;
			x_board_counter <= 8'b0;
			y_board_counter <= 8'b0;
			offset <= 8'b0;
			
			note1_bar <= note1_bar << 1;
			note2_bar <= note2_bar << 1;
			note3_bar <= note3_bar << 1;
			note4_bar <= note4_bar << 1;
			
			note1_bar[0] <= song_note1[818];
			note2_bar[0] <= song_note2[818];
			note3_bar[0] <= song_note3[818];
			note4_bar[0] <= song_note4[818];
			
			if(song_note1 == 819'b0 && song_note2 == 819'b0  && song_note3 == 819'b0  && song_note4 == 819'b0 )
				done <= 1'b0;
			else
				done <= 1'b1;
			
			if(shift_counter == 3'b100)
			begin
				song_note1 <= song_note1 << 1;
				song_note2 <= song_note2 << 1;
				song_note3 <= song_note3 << 1;
				song_note4 <= song_note4 << 1;
				shift_counter <= 3'b000;
			end
			else
				shift_counter <= shift_counter + 1'b1;
		
		end
		
		if(draw_board)
		begin
			updating <= 1'b1;
			colour_out <= 3'b111;
			offset <= 8'b0;
			
			if(x_board_counter < 8'd160 && line_counter == 4'b0000)
			begin
				x_coordinate <= x_board_counter;
				y_coordinate <= 8'd100;
				x_board_counter <= x_board_counter + 1'b1;
			end
			else if(x_board_counter < 8'd160 && line_counter == 4'b0001)
			begin
				x_coordinate <= x_board_counter;
				y_coordinate <= 8'd105;
				x_board_counter <= x_board_counter + 1'b1;
			end
			else if(y_board_counter < 8'd120 && line_counter == 4'b0010)
			begin
				x_coordinate <= 8'd0;
				y_coordinate <= y_board_counter;
				y_board_counter <= y_board_counter + 1'b1;
			end
			else if(y_board_counter < 8'd120 && line_counter == 4'b0011)
			begin
				x_coordinate <= 8'd40;
				y_coordinate <= y_board_counter;
				y_board_counter <= y_board_counter + 1'b1;
			end
			else if(y_board_counter < 8'd120 && line_counter == 4'b0100)
			begin
				x_coordinate <= 8'd80;
				y_coordinate <= y_board_counter;
				y_board_counter <= y_board_counter + 1'b1;
			end
			else if(y_board_counter < 8'd120 && line_counter == 4'b0101)
			begin
				x_coordinate <= 8'd120;
				y_coordinate <= y_board_counter;
				y_board_counter <= y_board_counter + 1'b1;
			end
			
			else if(y_board_counter < 8'd120 && line_counter == 4'b0111)
			begin
				x_coordinate <= 8'd159;
				y_coordinate <= y_board_counter;
				y_board_counter <= y_board_counter + 1'b1;
			end
			else
			begin
				line_counter <= line_counter + 1'b1;
				x_board_counter <= 8'b0;
				y_board_counter <= 8'b0;
				if(line_counter == 4'b0111)
				begin
					x_coordinate <= 8'b0;
					y_coordinate <= 8'b0;
					x_board_counter <= 8'b0;
					y_board_counter <= 8'b0;
					updating <= 1'b0;
					colour_out <= 3'b000;
				end
			end
			
		end
		
		if(draw_notes1)
		begin
		
			updating <= 1'b1;
			offset <= 8'd20;
			
			if(note1_bar[y_coordinate] == 1'b1)
				colour_out <= 3'b001;
			else if(y_coordinate == 8'd100 || y_coordinate == 8'd105)
				colour_out <= 3'b111;
			else
				colour_out <= 3'b000;
			
			
			if(counter < 3'b100)
			begin
				x_coordinate <= x_coordinate + 1'b1;
				counter <= counter + 1'b1;
			end
			else
			begin
				counter <= 3'b0;
				x_coordinate <= 8'b0;
				y_coordinate <= y_coordinate + 1'b1;
				if(y_coordinate == 8'b01111000)
				begin
					updating <= 1'b0;
					y_coordinate <= 8'b0;
					x_coordinate <= 8'b0;
				end
			
			end
			
		end
		
		
		if(draw_notes2)
		begin
			updating <= 1'b1;
			
			offset <= 8'd60;
			if(note2_bar[y_coordinate] == 1'b1)
				colour_out <= 3'b010;
			else if(y_coordinate == 8'd100 || y_coordinate == 8'd105)
				colour_out <= 3'b111;
			else
				colour_out <= 3'b000;
			
			
			if(counter < 3'b100)
			begin
				x_coordinate <= x_coordinate + 1'b1;
				counter <= counter + 1'b1;
			end
			else
			begin
				counter <= 3'b0;
				x_coordinate <= 8'b0;
				y_coordinate <= y_coordinate + 1'b1;
				if(y_coordinate == 8'b01111000)
				begin
					updating <= 1'b0;
					y_coordinate <= 8'b0;
					x_coordinate <= 8'b0;
				end
			
			end
			
		end
		
		if(draw_notes3)
		begin
			updating <= 1'b1;
			
			offset <= 8'd100;
			if(note3_bar[y_coordinate] == 1'b1)
				colour_out <= 3'b100;
			else if(y_coordinate == 8'd100 || y_coordinate == 8'd105)
				colour_out <= 3'b111;
			else
				colour_out <= 3'b000;
			
			
			if(counter < 3'b100)
			begin
				x_coordinate <= x_coordinate + 1'b1;
				counter <= counter + 1'b1;
			end
			else
			begin
				counter <= 3'b0;
				x_coordinate <= 8'b0;
				y_coordinate <= y_coordinate + 1'b1;
				if(y_coordinate == 8'b01111000)
				begin
					updating <= 1'b0;
					y_coordinate <= 8'b0;
					x_coordinate <= 8'b0;
				end
			
			end
			
		end
		
		if(draw_notes4)
		begin
			updating <= 1'b1;
			
			offset <= 8'd140;
			if(note4_bar[y_coordinate] == 1'b1)
				colour_out <= 3'b110;
			else if(y_coordinate == 8'd100 || y_coordinate == 8'd105)
				colour_out <= 3'b111;
			else
				colour_out <= 3'b000;
			
			
			if(counter < 3'b100)
			begin
				x_coordinate <= x_coordinate + 1'b1;
				counter <= counter + 1'b1;
			end
			else
			begin
				counter <= 3'b0;
				x_coordinate <= 8'b0;
				y_coordinate <= y_coordinate + 1'b1;
				if(y_coordinate == 8'b01111000)
				begin
					updating <= 1'b0;
					y_coordinate <= 8'b0;
					x_coordinate <= 8'b0;
				end
			
			end
			
		end
		
		if(check_notes)
		begin
		
			if(note1_bar[99] == 1'b0)
				next_note[0] <= 1'b1;
				
			if(note2_bar[99] == 1'b0)
				next_note[1] <= 1'b1;
			
			if(note3_bar[99] == 1'b0)
				next_note[2] <= 1'b1;
				
			if(note4_bar[99] == 1'b0)
				next_note[3] <= 1'b1;
		
		
			if(next_note[0] == 1'b1 && note1_bar[99] == 1'b1)
			begin
			
				if(note1_bar[95] == 1'b1)
					hold_note[0] <= 1'b1;
				else
					hold_note[0] <= 1'b0;
					
				next_note[0] <= 1'b0;
				
			end
			
			if(next_note[1] == 1'b1 && note2_bar[99] == 1'b1)
			begin
			
				if(note2_bar[95] == 1'b1)
					hold_note[1] <= 1'b1;
				else
					hold_note[1] <= 1'b0;
					
				next_note[1] <= 1'b0;
				
			end
			
			if(next_note[2] == 1'b1 && note3_bar[99] == 1'b1)
			begin
			
				if(note3_bar[95] == 1'b1)
					hold_note[2] <= 1'b1;
				else
					hold_note[2] <= 1'b0;
					
				next_note[2] <= 1'b0;
				
			end
			
			if(next_note[3] == 1'b1 && note4_bar[99] == 1'b1)
			begin
			
				if(note4_bar[95] == 1'b1)
					hold_note[3] <= 1'b1;
				else
					hold_note[3] <= 1'b0;
					
				next_note[3] <= 1'b0;
				
			end
				
			
		
		end
		
		if(playerEN)
		begin
		
			if(!keypress[3])
			begin
			
				if(note1_bar[100] == 1'b1 || note1_bar[101] == 1'b1 || note1_bar[102] == 1'b1 || note1_bar[103] == 1'b1)
				begin
				
					if(hold_note[0])
					begin
						note1_bar[10] <= 1'b0;
						temp_score1 <= temp_score1 + 1'b1;
					end
					else
					begin
						
						if(note1_bar[103] == 1'b1 && note1_bar[102] == 1'b1 && note1_bar[101] == 1'b1 && note1_bar[100] == 1'b1)
							temp_score1 <= temp_score1 + 4'd8;
						else if(note1_bar[100] == 1'b1 && note1_bar[101] == 1'b1 && note1_bar[102] == 1'b1)
							temp_score1 <= temp_score1 + 3'd4;
						else if(note1_bar[101] == 1'b1 && note1_bar[102] == 1'b1 && note1_bar[103] == 1'b1)
							temp_score1 <= temp_score1 + 3'd4;
						else if(note1_bar[101] == 1'b1 && note1_bar[100] == 1'b1)
							temp_score1 <= temp_score1 + 2'd2;
						else if(note1_bar[102] == 1'b1 && note1_bar[103] == 1'b1)
							temp_score1 <= temp_score1 + 2'd2;		
						else if(note1_bar[103] == 1'b1)
							temp_score1 <= temp_score1 + 1'd1;
						else if(note1_bar[100] == 1'b1)
							temp_score1 <= temp_score1 + 1'b1;
						
						
						if(note1_bar[99] == 1'b1);
						begin
							note1_bar[99] <= 1'b0;
							if(note1_bar[98] <= 1'b1)
							begin
								note1_bar[98] <= 1'b0;
								if(note1_bar[97] == 1'b1)
								begin
									note1_bar[97] <= 1'b0;
									if(note1_bar[96] == 1'b1)
										note1_bar[96] <= 1'b0;
								end
							end
						end
						
						note1_bar[100] <= 1'b0;
						note1_bar[101] <= 1'b0;
						note1_bar[102] <= 1'b0;
						note1_bar[103] <= 1'b0;
						note1_bar[104] <= 1'b0;
						note1_bar[105] <= 1'b0;
						note1_bar[106] <= 1'b0;
						note1_bar[107] <= 1'b0;
						
					end
				
					colour_out <= 3'b000;
					
				end
				
				
				
			end
			
			if(!keypress[2])
			begin
				if(note2_bar[100] == 1'b1 || note2_bar[101] == 1'b1 || note2_bar[102] == 1'b1 || note2_bar[103] == 1'b1)
				begin
				
					if(hold_note[1])
					begin
						note2_bar[103] <= 1'b0;
						temp_score2 <= temp_score2 + 1'b1;
					end
					else
					begin
						
						if(note2_bar[103] == 1'b1 && note2_bar[102] == 1'b1 && note2_bar[101] == 1'b1 && note2_bar[100] == 1'b1)
							temp_score2 <= temp_score2 + 4'd8;
						else if(note2_bar[100] == 1'b1 && note2_bar[101] == 1'b1 && note2_bar[102] == 1'b1)
							temp_score2 <= temp_score2 + 3'd4;
						else if(note2_bar[101] == 1'b1 && note2_bar[102] == 1'b1 && note2_bar[103] == 1'b1)
							temp_score2 <= temp_score2 + 3'd4;
						else if(note2_bar[101] == 1'b1 && note2_bar[100] == 1'b1)
							temp_score2 <= temp_score2 + 2'd2;
						else if(note2_bar[102] == 1'b1 && note2_bar[103] == 1'b1)
							temp_score2 <= temp_score2 + 2'd2;		
						else if(note2_bar[103] == 1'b1)
							temp_score2 <= temp_score2 + 1'd1;
						else if(note2_bar[100] == 1'b1)
							temp_score2 <= temp_score2 + 1'b1;
						
						
						if(note2_bar[99] == 1'b1);
						begin
							note2_bar[99] <= 1'b0;
							if(note2_bar[98] <= 1'b1)
							begin
								note2_bar[98] <= 1'b0;
								if(note2_bar[97] == 1'b1)
								begin
									note2_bar[97] <= 1'b0;
									if(note2_bar[96] == 1'b1)
										note2_bar[96] <= 1'b0;
								end
							end
						end
						
						note2_bar[100] <= 1'b0;
						note2_bar[101] <= 1'b0;
						note2_bar[102] <= 1'b0;
						note2_bar[103] <= 1'b0;
						note2_bar[104] <= 1'b0;
						note2_bar[105] <= 1'b0;
						note2_bar[106] <= 1'b0;
						note2_bar[107] <= 1'b0;
						
					end
				
					colour_out <= 3'b000;
					
				end
			end
			
			if(!keypress[1])
			begin
				if(note3_bar[100] == 1'b1 || note3_bar[101] == 1'b1 || note3_bar[102] == 1'b1 || note3_bar[103] == 1'b1)
				begin
				
					if(hold_note[2])
					begin
						note3_bar[103] <= 1'b0;
						temp_score3 <= temp_score3 + 1'b1;
					end
					else
					begin
						
						if(note3_bar[103] == 1'b1 && note3_bar[102] == 1'b1 && note3_bar[101] == 1'b1 && note3_bar[100] == 1'b1)
							temp_score3 <= temp_score3 + 4'd8;
						else if(note3_bar[100] == 1'b1 && note3_bar[101] == 1'b1 && note3_bar[102] == 1'b1)
							temp_score3 <= temp_score3 + 3'd4;
						else if(note3_bar[101] == 1'b1 && note3_bar[102] == 1'b1 && note3_bar[103] == 1'b1)
							temp_score3 <= temp_score3 + 3'd4;
						else if(note3_bar[101] == 1'b1 && note3_bar[100] == 1'b1)
							temp_score3 <= temp_score3 + 2'd2;
						else if(note3_bar[102] == 1'b1 && note3_bar[103] == 1'b1)
							temp_score3 <= temp_score3 + 2'd2;		
						else if(note3_bar[103] == 1'b1)
							temp_score3 <= temp_score3 + 1'd1;
						else if(note3_bar[100] == 1'b1)
							temp_score3 <= temp_score3 + 1'b1;
						
						
						if(note3_bar[99] == 1'b1);
						begin
							note3_bar[99] <= 1'b0;
							if(note3_bar[98] <= 1'b1)
							begin
								note3_bar[98] <= 1'b0;
								if(note3_bar[97] == 1'b1)
								begin
									note3_bar[97] <= 1'b0;
									if(note3_bar[96] == 1'b1)
										note3_bar[96] <= 1'b0;
								end
							end
						end
						
						note3_bar[100] <= 1'b0;
						note3_bar[101] <= 1'b0;
						note3_bar[102] <= 1'b0;
						note3_bar[103] <= 1'b0;
						note3_bar[104] <= 1'b0;
						note3_bar[105] <= 1'b0;
						note3_bar[106] <= 1'b0;
						note3_bar[107] <= 1'b0;
						
					end
				
					colour_out <= 3'b000;
					
				end
			end
			
			if(!keypress[0])
			begin
				if(note4_bar[100] == 1'b1 || note4_bar[101] == 1'b1 || note4_bar[102] == 1'b1 || note4_bar[103] == 1'b1)
				begin
				
					if(hold_note[3])
					begin
						note4_bar[103] <= 1'b0;
						temp_score4 <= temp_score4 + 1'b1;
					end
					else
					begin
						
						if(note4_bar[103] == 1'b1 && note4_bar[102] == 1'b1 && note4_bar[101] == 1'b1 && note4_bar[100] == 1'b1)
							temp_score4 <= temp_score4 + 4'd8;
						else if(note4_bar[100] == 1'b1 && note4_bar[101] == 1'b1 && note4_bar[102] == 1'b1)
							temp_score4 <= temp_score4 + 3'd4;
						else if(note4_bar[101] == 1'b1 && note4_bar[102] == 1'b1 && note4_bar[103] == 1'b1)
							temp_score4 <= temp_score4 + 3'd4;
						else if(note4_bar[101] == 1'b1 && note4_bar[100] == 1'b1)
							temp_score4 <= temp_score4 + 2'd2;
						else if(note4_bar[102] == 1'b1 && note4_bar[103] == 1'b1)
							temp_score4 <= temp_score4 + 2'd2;		
						else if(note4_bar[103] == 1'b1)
							temp_score4 <= temp_score4 + 1'd1;
						else if(note4_bar[100] == 1'b1)
							temp_score4 <= temp_score4 + 1'b1;
						
						
						if(note4_bar[99] == 1'b1);
						begin
							note4_bar[99] <= 1'b0;
							if(note4_bar[98] <= 1'b1)
							begin
								note4_bar[98] <= 1'b0;
								if(note4_bar[97] == 1'b1)
								begin
									note4_bar[97] <= 1'b0;
									if(note4_bar[96] == 1'b1)
										note4_bar[96] <= 1'b0;
								end
							end
						end
						
						note4_bar[100] <= 1'b0;
						note4_bar[101] <= 1'b0;
						note4_bar[102] <= 1'b0;
						note4_bar[103] <= 1'b0;
						note4_bar[104] <= 1'b0;
						note4_bar[105] <= 1'b0;
						note4_bar[106] <= 1'b0;
						note4_bar[107] <= 1'b0;
						
					end
				
					colour_out <= 3'b000;
					
				end
			end
		
		end
		
		score <= temp_score1 + temp_score2 + temp_score3 + temp_score4;
		x_out <= x_coordinate + offset;
		y_out <= y_coordinate;
		
	end
	
	
endmodule
